module dec_counter(output reg [3:0]count,input clk,reset);
  //????
  always@(posedge clk)begin
    if(reset)
      count<=4'b0;
    else if(count==4'b1010)
      //????????????0~9??0~10??????9
      //???10????4'b1010
      count<=4'b0;
    else
      count<=count+1'b1;
  end
endmodule
